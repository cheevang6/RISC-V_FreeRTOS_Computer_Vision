module svTest();

enum {one,two,three} number;

endmodule