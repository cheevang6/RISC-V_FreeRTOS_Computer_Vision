//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Fri Dec  4 17:33:41 2020
// Version: v12.3 12.800.0.16
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// sccb_design
module sccb_design(
    // Inputs
    xclk,
    // Outputs
    sio_c,
    // Inouts
    sio_d
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input  xclk;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output sio_c;
//--------------------------------------------------------------------
// Inout
//--------------------------------------------------------------------
inout  sio_d;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire   sio_c_net_0;
wire   sio_d;
wire   xclk;
wire   sio_c_net_1;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire   VCC_net;
wire   [7:0]data_in_const_net_0;
wire   [7:0]addr_id_const_net_0;
wire   [7:0]addr_reg_const_net_0;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign VCC_net              = 1'b1;
assign data_in_const_net_0  = 8'h00;
assign addr_id_const_net_0  = 8'h00;
assign addr_reg_const_net_0 = 8'h00;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign sio_c_net_1 = sio_c_net_0;
assign sio_c       = sio_c_net_1;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------SCCB_CTRL
SCCB_CTRL SCCB_CTRL_0(
        // Inputs
        .XCLK     ( xclk ),
        .RST_N    ( VCC_net ),
        .RW       ( VCC_net ),
        .data_in  ( data_in_const_net_0 ),
        .addr_id  ( addr_id_const_net_0 ),
        .addr_reg ( addr_reg_const_net_0 ),
        // Outputs
        .SIO_C    ( sio_c_net_0 ),
        .data_out (  ),
        // Inouts
        .SIO_D    ( sio_d ) 
        );


endmodule
